../../tb_tcdm_interconnect/hdl/tb_pkg.sv