// Copyright 2021 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

`include "axi/assign.svh"
`include "common_cells/registers.svh"

module mempool_system
  import mempool_pkg::*;
#(
  // TCDM
  parameter addr_t       TCDMBaseAddr  = 32'h0000_0000,
  // Boot address
  parameter addr_t       BootAddr      = 32'h0000_0000
) (
  input logic                clk_i,
  input logic                rst_ni,

  input  logic               fetch_en_i,
  output logic               eoc_valid_o,
  output logic               busy_o,

  output axi_system_req_t    mst_req_o,
  input  axi_system_resp_t   mst_resp_i,

  input  axi_system_req_t    slv_req_i,
  output axi_system_resp_t   slv_resp_o
);

  import axi_pkg::xbar_cfg_t;
  import axi_pkg::xbar_rule_32_t;

  /*********
   *  AXI  *
   *********/

  // Overview of AXI buses with SRAM L2
  //
  //      mst_demux
  //        / |
  //       /  | soc  +----------+ periph  +---------+
  //      |  0|=====>| soc_xbar |========>| periph  |
  //  mst |   |      +----------+         +---------+
  // ====>|   |
  //      |   | l2   +----------+  mem    +---------+ bank  +--------+
  //      |  1|=====>| axi2mem  |-------->| l2_xbar |------>| l2_mem |
  //       \  |      +----------+         +---------+       +--------+
  //        \_|
  //                  == axi ==>          -- tcdm -->
  //
  // Overview of AXI buses with DRAM L2
  //
  //      mst_demux
  //        / |
  //       /  | soc  +----------+ periph  +---------+
  //      |  0|=====>| soc_xbar |========>| periph  |
  //  mst |   |      +----------+         +---------+
  // ====>|   |
  //      |   | l2   +----------+  mem_one_port  +--------------+
  //      |  1|=====>| AXI_Mux  |===============>| AXI Port Out |
  //       \  |      +----------+                +--------------+
  //        \_|
  //                  == axi ==>

  localparam NumAXISlaves  = 3; // control regs, bootrom and the external mst ports
  localparam NumSoCRules   = NumAXISlaves - 1;

  typedef enum logic [$clog2(NumAXISlaves) - 1:0] {
    Peripherals,
    Bootrom,
    External
  } axi_soc_xbar_slave_target;

  typedef enum logic {
    SoCXBar = 0,
    L2Memory = 1
  } axi_mst_demux_slave_target;

  axi_tile_req_t    [NumSystemXbarMasters-1:0] axi_mst_req;
  axi_tile_resp_t   [NumSystemXbarMasters-1:0] axi_mst_resp;
  axi_tile_req_t    [NumSystemXbarMasters-1:0] axi_cluster_req;
  axi_tile_req_t    [NumSystemXbarMasters-1:0] axi_l2_req;
  axi_tile_resp_t   [NumSystemXbarMasters-1:0] axi_l2_resp;
  axi_tile_req_t    [NumSystemXbarMasters-1:0] axi_soc_req;
  axi_tile_resp_t   [NumSystemXbarMasters-1:0] axi_soc_resp;
  axi_system_req_t  [NumAXISlaves-1:0]  axi_periph_req;
  axi_system_resp_t [NumAXISlaves-1:0]  axi_periph_resp;

  logic             [NumClusters-1:0][NumCores-1:0]      wake_up;
  logic             [NumClusters-1:0]                    eoc_valid;
  ro_cache_ctrl_t   [NumClusters-1:0]                    ro_cache_ctrl;
  dma_req_t  [NumClusters-1:0]dma_req;
  logic      [NumClusters-1:0]dma_req_valid;
  logic      [NumClusters-1:0]dma_req_ready;
  dma_meta_t [NumClusters-1:0]dma_meta;
  logic      [NumClusters-1:0][1-1:0] dma_id;

  localparam xbar_cfg_t MstDemuxCfg = '{
    NoSlvPorts         : 1, // Each master has a private demux
    NoMstPorts         : 2, // going to either the xbar or L2
    MaxMstTrans        : 4,
    MaxSlvTrans        : 4,
    FallThrough        : 1'b0,
    LatencyMode        : axi_pkg::NO_LATENCY,
    PipelineStages     : 0,
    AxiIdWidthSlvPorts : AxiTileIdWidth,
    AxiIdUsedSlvPorts  : AxiTileIdWidth,
    UniqueIds          : 0,
    AxiAddrWidth       : AddrWidth,
    AxiDataWidth       : AxiDataWidth,
    NoAddrRules        : 1
  };

  localparam xbar_cfg_t SoCXBarCfg = '{
    NoSlvPorts         : NumSystemXbarMasters,
    NoMstPorts         : NumAXISlaves,
    MaxMstTrans        : 4,
    MaxSlvTrans        : 4,
    FallThrough        : 1'b0,
    LatencyMode        : axi_pkg::CUT_MST_PORTS,
    PipelineStages     : 0,
    AxiIdWidthSlvPorts : AxiTileIdWidth,
    AxiIdUsedSlvPorts  : AxiTileIdWidth,
    UniqueIds          : 0,
    AxiAddrWidth       : AddrWidth,
    AxiDataWidth       : AxiDataWidth,
    NoAddrRules        : NumSoCRules
  };

  /*********************
   *  MemPool Cluster  *
   ********************/
  assign eoc_valid_o = eoc_valid[0];
  for(genvar i = 0; i < NumClusters; i++) begin: gen_clusters
    mempool_cluster #(
      .TCDMBaseAddr(TCDMBaseAddr),
      .BootAddr    (BootAddr    )
    ) i_mempool_cluster (
      .clk_i          (clk_i                          ),
      .rst_ni         (rst_ni                         ),
      .cluster_id_i   (i                              ),
      .wake_up_i      (wake_up[i]                     ),
      .testmode_i     (1'b0                           ),
      .scan_enable_i  (1'b0                           ),
      .scan_data_i    (1'b0                           ),
      .scan_data_o    (/* Unused */                   ),
      .ro_cache_ctrl_i(ro_cache_ctrl[i]                  ),
      .dma_req_i      (dma_req[i]                        ),
      .dma_req_valid_i(dma_req_valid[i]                  ),
      .dma_req_ready_o(dma_req_ready[i]                  ),
      .dma_meta_o     (dma_meta[i]                       ),
      .axi_mst_req_o  (axi_cluster_req[i*NumClusterAXIMasters +: NumClusterAXIMasters] ),
      .axi_mst_resp_i (axi_mst_resp[i*NumClusterAXIMasters +: NumClusterAXIMasters])
    );

    for(genvar j = 0; j < NumClusterAXIMasters; j++) begin: gen_axi_assignment
      // address_write
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.id = axi_cluster_req[i*NumClusterAXIMasters+j].aw.id;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.addr = axi_cluster_req[i*NumClusterAXIMasters+j].aw.addr;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.len = axi_cluster_req[i*NumClusterAXIMasters+j].aw.len;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.size = axi_cluster_req[i*NumClusterAXIMasters+j].aw.size;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.burst = axi_cluster_req[i*NumClusterAXIMasters+j].aw.burst;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.lock = axi_cluster_req[i*NumClusterAXIMasters+j].aw.lock;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.cache = axi_cluster_req[i*NumClusterAXIMasters+j].aw.cache;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.prot = axi_cluster_req[i*NumClusterAXIMasters+j].aw.prot;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.qos = axi_cluster_req[i*NumClusterAXIMasters+j].aw.qos;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.region = axi_cluster_req[i*NumClusterAXIMasters+j].aw.region;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.atop = axi_cluster_req[i*NumClusterAXIMasters+j].aw.atop;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw.user = i;
      // address_read
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.id = axi_cluster_req[i*NumClusterAXIMasters+j].ar.id;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.addr = axi_cluster_req[i*NumClusterAXIMasters+j].ar.addr;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.len = axi_cluster_req[i*NumClusterAXIMasters+j].ar.len;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.size = axi_cluster_req[i*NumClusterAXIMasters+j].ar.size;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.burst = axi_cluster_req[i*NumClusterAXIMasters+j].ar.burst;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.lock = axi_cluster_req[i*NumClusterAXIMasters+j].ar.lock;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.cache = axi_cluster_req[i*NumClusterAXIMasters+j].ar.cache;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.prot = axi_cluster_req[i*NumClusterAXIMasters+j].ar.prot;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.qos = axi_cluster_req[i*NumClusterAXIMasters+j].ar.qos;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.region = axi_cluster_req[i*NumClusterAXIMasters+j].ar.region;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar.user = i;
      assign axi_mst_req[i*NumClusterAXIMasters+j].aw_valid = axi_cluster_req[i*NumClusterAXIMasters+j].aw_valid;
      assign axi_mst_req[i*NumClusterAXIMasters+j].w = axi_cluster_req[i*NumClusterAXIMasters+j].w;
      assign axi_mst_req[i*NumClusterAXIMasters+j].w_valid = axi_cluster_req[i*NumClusterAXIMasters+j].w_valid;
      assign axi_mst_req[i*NumClusterAXIMasters+j].b_ready = axi_cluster_req[i*NumClusterAXIMasters+j].b_ready;
      assign axi_mst_req[i*NumClusterAXIMasters+j].ar_valid = axi_cluster_req[i*NumClusterAXIMasters+j].ar_valid;
      assign axi_mst_req[i*NumClusterAXIMasters+j].r_ready = axi_cluster_req[i*NumClusterAXIMasters+j].r_ready;
    end

  end

  /**********************
   *  AXI Interconnect  *
   **********************/

  localparam addr_t PeripheralsBaseAddr   = 32'h4000_0000;
  localparam addr_t PeripheralsEndAddr    = 32'h4002_0000;
  localparam addr_t L2MemoryBaseAddr      = `ifdef L2_BASE `L2_BASE `else 32'h8000_0000 `endif;
  localparam addr_t L2MemoryEndAddr       = L2MemoryBaseAddr + L2Size;
  localparam addr_t BootromBaseAddr       = 32'hA000_0000;
  localparam addr_t BootromEndAddr        = 32'hA000_FFFF;

  xbar_rule_32_t [            0:0]  mst_demux_rules;
  xbar_rule_32_t [NumSoCRules-1:0] soc_xbar_rules;
  assign mst_demux_rules = '{
    '{idx: L2Memory, start_addr: L2MemoryBaseAddr, end_addr: L2MemoryEndAddr}
  };
  assign soc_xbar_rules = '{
    '{idx: Peripherals, start_addr: PeripheralsBaseAddr, end_addr: PeripheralsEndAddr},
    '{idx: Bootrom, start_addr: BootromBaseAddr, end_addr: BootromEndAddr}
  };

  for (genvar i = 0; i < NumSystemXbarMasters; i++) begin : gen_mst_demux
    axi_xbar #(
      .Cfg          (MstDemuxCfg      ),
      .slv_aw_chan_t(axi_tile_aw_t    ),
      .mst_aw_chan_t(axi_tile_aw_t    ),
      .w_chan_t     (axi_tile_w_t     ),
      .slv_b_chan_t (axi_tile_b_t     ),
      .mst_b_chan_t (axi_tile_b_t     ),
      .slv_ar_chan_t(axi_tile_ar_t    ),
      .mst_ar_chan_t(axi_tile_ar_t    ),
      .slv_r_chan_t (axi_tile_r_t     ),
      .mst_r_chan_t (axi_tile_r_t     ),
      .slv_req_t    (axi_tile_req_t   ),
      .slv_resp_t   (axi_tile_resp_t  ),
      .mst_req_t    (axi_tile_req_t   ),
      .mst_resp_t   (axi_tile_resp_t  ),
      .rule_t       (xbar_rule_32_t   )
    ) i_mst_demux (
      .clk_i                (clk_i                           ),
      .rst_ni               (rst_ni                          ),
      .test_i               (1'b0                            ),
      .slv_ports_req_i      (axi_mst_req[i]                  ),
      .slv_ports_resp_o     (axi_mst_resp[i]                 ),
      .mst_ports_req_o      ({axi_l2_req[i] ,axi_soc_req[i] }),
      .mst_ports_resp_i     ({axi_l2_resp[i],axi_soc_resp[i]}),
      .addr_map_i           (mst_demux_rules                 ),
      .en_default_mst_port_i(1'b1                            ),
      .default_mst_port_i   (SoCXBar                         )
    );
  end

  axi_xbar #(
    .Cfg          (SoCXBarCfg       ),
    .slv_aw_chan_t(axi_tile_aw_t    ),
    .mst_aw_chan_t(axi_system_aw_t  ),
    .w_chan_t     (axi_tile_w_t     ),
    .slv_b_chan_t (axi_tile_b_t     ),
    .mst_b_chan_t (axi_system_b_t   ),
    .slv_ar_chan_t(axi_tile_ar_t    ),
    .mst_ar_chan_t(axi_system_ar_t  ),
    .slv_r_chan_t (axi_tile_r_t     ),
    .mst_r_chan_t (axi_system_r_t   ),
    .slv_req_t    (axi_tile_req_t   ),
    .slv_resp_t   (axi_tile_resp_t  ),
    .mst_req_t    (axi_system_req_t ),
    .mst_resp_t   (axi_system_resp_t),
    .rule_t       (xbar_rule_32_t   )
  ) i_soc_xbar (
    .clk_i                (clk_i                    ),
    .rst_ni               (rst_ni                   ),
    .test_i               (1'b0                     ),
    .slv_ports_req_i      (axi_soc_req              ),
    .slv_ports_resp_o     (axi_soc_resp             ),
    .mst_ports_req_o      (axi_periph_req           ),
    .mst_ports_resp_i     (axi_periph_resp          ),
    .addr_map_i           (soc_xbar_rules           ),
    .en_default_mst_port_i({NumSystemXbarMasters{1'b1}}    ), // default all slave ports to master port External
    .default_mst_port_i   ({NumSystemXbarMasters{External}})
  );

`ifndef DRAM

  /*************
   *  L2 SRAM  *
   *************/

  localparam int unsigned NumAXIMastersLog2 = NumSystemXbarMasters == 1 ? 1 : $clog2(NumSystemXbarMasters);
  typedef logic [L2AddrWidth-1:0] l2_mem_addr_t;
  typedef logic [L2BankAddrWidth-1:0] l2_bank_addr_t;
  typedef logic [NumAXIMastersLog2-1:0] bank_ini_t;
  // Axi2Mems to l2_xbar
  logic         [NumSystemXbarMasters-1:0] mem_req;
  logic         [NumSystemXbarMasters-1:0] mem_gnt;
  logic         [NumSystemXbarMasters-1:0] mem_rvalid;
  addr_t        [NumSystemXbarMasters-1:0] mem_addr_full;
  l2_mem_addr_t [NumSystemXbarMasters-1:0] mem_addr;
  axi_data_t    [NumSystemXbarMasters-1:0] mem_wdata;
  axi_strb_t    [NumSystemXbarMasters-1:0] mem_strb;
  logic         [NumSystemXbarMasters-1:0] mem_we;
  axi_data_t    [NumSystemXbarMasters-1:0] mem_rdata;
  // l2_xbar to banks
  logic          [NumL2Banks-1:0] bank_req;
  logic          [NumL2Banks-1:0] bank_gnt;
  logic          [NumL2Banks-1:0] bank_rvalid;
  l2_bank_addr_t [NumL2Banks-1:0] bank_addr;
  bank_ini_t     [NumL2Banks-1:0] bank_ini_d, bank_ini_q;
  axi_data_t     [NumL2Banks-1:0] bank_wdata;
  axi_strb_t     [NumL2Banks-1:0] bank_strb;
  logic          [NumL2Banks-1:0] bank_we;
  axi_data_t     [NumL2Banks-1:0] bank_rdata;

  for (genvar i = 0; i < NumSystemXbarMasters; i++) begin : gen_l2_adapters
    axi2mem #(
      .axi_req_t (axi_tile_req_t ),
      .axi_resp_t(axi_tile_resp_t),
      .AddrWidth (L2AddrWidth    ),
      .DataWidth (AxiDataWidth   ),
      .IdWidth   (AxiTileIdWidth ),
      .NumBanks  (1              ),
      .BufDepth  (3              )
    ) i_axi2mem (
      .clk_i       (clk_i         ),
      .rst_ni      (rst_ni        ),
      .busy_o      (/*unsused*/   ),
      .axi_req_i   (axi_l2_req[i] ),
      .axi_resp_o  (axi_l2_resp[i]),
      .mem_req_o   (mem_req[i]    ),
      .mem_gnt_i   (mem_gnt[i]    ),
      .mem_addr_o  (mem_addr[i]   ),
      .mem_wdata_o (mem_wdata[i]  ),
      .mem_strb_o  (mem_strb[i]   ),
      .mem_atop_o  (/*unused*/    ),
      .mem_we_o    (mem_we[i]     ),
      .mem_rvalid_i(mem_rvalid[i] ),
      .mem_rdata_i (mem_rdata[i]  )
    );
  end

  variable_latency_interconnect #(
    .NumIn            (NumSystemXbarMasters  ),
    .NumOut           (NumL2Banks     ),
    .AddrWidth        (L2AddrWidth    ),
    .DataWidth        (L2BankWidth    ),
    .BeWidth          (L2BankBeWidth  ),
    .AddrMemWidth     (L2BankAddrWidth),
    .AxiVldRdy        (1'b1           ),
    .SpillRegisterReq (64'b1          ),
    .SpillRegisterResp(64'b1          )
  ) i_l2_xbar (
    .clk_i          (clk_i      ),
    .rst_ni         (rst_ni     ),
    // master side
    .req_valid_i    (mem_req    ),
    .req_ready_o    (mem_gnt    ),
    .req_tgt_addr_i (mem_addr   ),
    .req_wen_i      (mem_we     ),
    .req_wdata_i    (mem_wdata  ),
    .req_be_i       (mem_strb   ),
    .resp_valid_o   (mem_rvalid ),
    .resp_ready_i   ('1         ),
    .resp_rdata_o   (mem_rdata  ),
    // slave side
    .req_valid_o    (bank_req   ),
    .req_ready_i    ('1         ),
    .req_ini_addr_o (bank_ini_d ),
    .req_tgt_addr_o (bank_addr  ),
    .req_wen_o      (bank_we    ),
    .req_wdata_o    (bank_wdata ),
    .req_be_o       (bank_strb  ),
    .resp_valid_i   (bank_rvalid),
    .resp_ready_o   (/*unused*/ ), // This only works because resp_ready_i = 1
    .resp_ini_addr_i(bank_ini_q ),
    .resp_rdata_i   (bank_rdata )
  );

  `FF(bank_rvalid, bank_req, 1'b0, clk_i, rst_ni)
  `FF(bank_ini_q, bank_ini_d, 1'b0, clk_i, rst_ni)

  // The initialization at reset is not supported by Verilator. Therefore, we disable the SimInit at
  // reset for Verilator. Since our preloading through the SystemVerilog testbench requires the
  // SimInit value to be assigned at reset, we use the "custom" string to invoke the initialization
  // without setting the memory to known values like "ones" or "zeros".
  localparam L2SimInit = `ifdef VERILATOR "none" `else "custom" `endif;
  for (genvar i = 0; i < NumL2Banks; i++) begin : gen_l2_banks
    tc_sram #(
      .DataWidth(L2BankWidth   ),
      .NumWords (L2BankNumWords),
      .NumPorts (1             ),
      .SimInit  (L2SimInit     )
    ) l2_mem (
      .clk_i  (clk_i        ),
      .rst_ni (rst_ni       ),
      .req_i  (bank_req[i]  ),
      .we_i   (bank_we[i]   ),
      .addr_i (bank_addr[i] ),
      .wdata_i(bank_wdata[i]),
      .be_i   (bank_strb[i] ),
      .rdata_o(bank_rdata[i])
    );
  end

`else

  /*************
   *  L2 DRAM  *
   *************/

  // AXI xbar to form one port to DRAM
  localparam NumDramRules = NumDrams;

  xbar_rule_32_t    [NumDramRules-1:0] dram_xbar_rules;
  axi_system_req_t  [NumDrams-1:0]     dram_req_interleaved;
  axi_system_req_t  [NumDrams-1:0]     dram_req;
  axi_system_resp_t [NumDrams-1:0]     dram_resp;

  // AXI brust splitter for DRAM interleaving
  axi_tile_req_t  [NumSystemXbarMasters-1:0] axi_l2_req_splitted;
  axi_tile_resp_t [NumSystemXbarMasters-1:0] axi_l2_resp_splitted;
  axi_tile_req_t  [NumSystemXbarMasters-1:0] axi_l2_req_interleaved;

  generate
    if (DmaBrustLen > Interleave) begin : gen_axi_splitter
      for (genvar i = 0; unsigned'(i) < NumSystemXbarMasters; i++) begin: brust_splitter
        axi_burst_splitter #(
          .MaxReadTxns (16             ),
          .MaxWriteTxns(16             ),
          .AddrWidth   (AddrWidth      ),
          .DataWidth   (AxiDataWidth   ),
          .IdWidth     (AxiTileIdWidth ),
          .UserWidth   (1              ),
          .axi_req_t   (axi_tile_req_t ),
          .axi_resp_t  (axi_tile_resp_t)
        ) i_axi_burst_splitter (
          .clk_i     (clk_i                  ),
          .rst_ni    (rst_ni                 ),
          .slv_req_i (axi_l2_req[i]          ),
          .slv_resp_o(axi_l2_resp[i]         ),
          .mst_req_o (axi_l2_req_splitted[i] ),
          .mst_resp_i(axi_l2_resp_splitted[i])
        );
      end: brust_splitter
    end else begin : splitter_bypass
      // Do not need a splitter
      assign axi_l2_req_splitted  = axi_l2_req;
      assign axi_l2_resp          = axi_l2_resp_splitted;
    end: splitter_bypass
  endgenerate

  localparam int unsigned ConstantBits = $clog2(L2BankBeWidth * Interleave);
  localparam int unsigned ScrambleBits = (NumDrams == 1) ? 1 : $clog2(NumDrams);
  localparam int unsigned ReminderBits = AddrWidth - ScrambleBits - ConstantBits;
  // req.aw scrambling
  logic [NumSystemXbarMasters-1:0][ConstantBits-1:0] aw_const;
  logic [NumSystemXbarMasters-1:0][ScrambleBits-1:0] aw_scramble;
  logic [NumSystemXbarMasters-1:0][ReminderBits-1:0] aw_reminder;
  logic [NumSystemXbarMasters-1:0][AddrWidth-1   :0] aw_scramble_addr;
  // req.ar scrambling
  logic [NumSystemXbarMasters-1:0][ConstantBits-1:0] ar_const;
  logic [NumSystemXbarMasters-1:0][ScrambleBits-1:0] ar_scramble;
  logic [NumSystemXbarMasters-1:0][ReminderBits-1:0] ar_reminder;
  logic [NumSystemXbarMasters-1:0][AddrWidth-1   :0] ar_scramble_addr;

  for (genvar i = 0; unsigned'(i) < NumSystemXbarMasters; i++) begin: gen_dram_scrambler
    assign aw_const[i]         = axi_l2_req_splitted[i].aw.addr[ConstantBits-1 : 0];
    assign aw_scramble[i]      = axi_l2_req_splitted[i].aw.addr[ScrambleBits+ConstantBits-1 : ConstantBits];
    assign aw_reminder[i]      = axi_l2_req_splitted[i].aw.addr[AddrWidth-1 : ScrambleBits+ConstantBits];
    assign aw_scramble_addr[i] = {aw_scramble[i], aw_reminder[i], aw_const[i]};

    assign ar_const[i]         = axi_l2_req_splitted[i].ar.addr[ConstantBits-1 : 0];
    assign ar_scramble[i]      = axi_l2_req_splitted[i].ar.addr[ScrambleBits+ConstantBits-1 : ConstantBits];
    assign ar_reminder[i]      = axi_l2_req_splitted[i].ar.addr[AddrWidth-1 : ScrambleBits+ConstantBits];
    assign ar_scramble_addr[i] = {ar_scramble[i], ar_reminder[i], ar_const[i]};

    // Scrambled AXI req assignment
    always_comb begin
      axi_l2_req_interleaved[i]         = axi_l2_req_splitted[i];
      axi_l2_req_interleaved[i].aw.addr = aw_scramble_addr[i];
      axi_l2_req_interleaved[i].ar.addr = ar_scramble_addr[i];
    end
  end: gen_dram_scrambler

  // DRAM Xbar rules
  for (genvar i = 0; unsigned'(i) < NumDramRules; i++) begin: gen_dram_xbar_rules
    logic [AddrWidth-1:0] start_dram_addr;
    logic [AddrWidth-1:0] end_dram_addr;
    assign start_dram_addr    = {{ScrambleBits{i}}, 1'b1, {AddrWidth-ScrambleBits-1{1'b0}}};
    assign end_dram_addr      = {{ScrambleBits{i}}, 1'b1, {AddrWidth-ScrambleBits-1{1'b1}}};
    assign dram_xbar_rules[i] = '{idx: i, start_addr: start_dram_addr, end_addr: end_dram_addr};
  end: gen_dram_xbar_rules

  // AXI Crossbar
  localparam xbar_cfg_t DRAMXBarCfg = '{
    NoSlvPorts         : NumSystemXbarMasters,
    NoMstPorts         : NumDrams,
    MaxMstTrans        : 16,
    MaxSlvTrans        : 16,
    FallThrough        : 16,
    LatencyMode        : axi_pkg::CUT_MST_PORTS,
    AxiIdWidthSlvPorts : AxiTileIdWidth,
    AxiIdUsedSlvPorts  : AxiTileIdWidth,
    UniqueIds          : 0,
    AxiAddrWidth       : AddrWidth,
    AxiDataWidth       : AxiDataWidth,
    NoAddrRules        : NumDramRules
  };

  axi_xbar #(
    .Cfg          (DRAMXBarCfg      ),
    .slv_aw_chan_t(axi_tile_aw_t    ),
    .mst_aw_chan_t(axi_system_aw_t  ),
    .w_chan_t     (axi_system_w_t   ),
    .slv_b_chan_t (axi_tile_b_t     ),
    .mst_b_chan_t (axi_system_b_t   ),
    .slv_ar_chan_t(axi_tile_ar_t    ),
    .mst_ar_chan_t(axi_system_ar_t  ),
    .slv_r_chan_t (axi_tile_r_t     ),
    .mst_r_chan_t (axi_system_r_t   ),
    .slv_req_t    (axi_tile_req_t   ),
    .slv_resp_t   (axi_tile_resp_t  ),
    .mst_req_t    (axi_system_req_t ),
    .mst_resp_t   (axi_system_resp_t),
    .rule_t       (xbar_rule_32_t   )
  ) i_dram_xbar (
    .clk_i                (clk_i                 ),
    .rst_ni               (rst_ni                ),
    .test_i               (1'b0                  ),
    .slv_ports_req_i      (axi_l2_req_interleaved),
    .slv_ports_resp_o     (axi_l2_resp_splitted  ),
    .mst_ports_req_o      (dram_req_interleaved  ),
    .mst_ports_resp_i     (dram_resp             ),
    .addr_map_i           (dram_xbar_rules       ),
    .en_default_mst_port_i({NumSystemXbarMasters{1'b1}} ),
    .default_mst_port_i   ('0                    )
  );

  // Scrambled Addr reset, and detect base address before go to DRAM
  for (genvar i = 0; unsigned'(i) < NumDrams; i++) begin: gen_dram_scrambler_reset
    // req.aw scrambling
    logic [ConstantBits-1:0] aw_const;
    logic [ScrambleBits-1:0] aw_scramble;
    logic [ReminderBits-1:0] aw_reminder;
    logic [AddrWidth-1   :0] aw_scramble_addr_reset;
    assign aw_scramble = dram_req_interleaved[i].aw.addr[AddrWidth-1 : AddrWidth-ScrambleBits];
    assign aw_reminder = dram_req_interleaved[i].aw.addr[AddrWidth-ScrambleBits-1 : ConstantBits] - L2MemoryBaseAddr[AddrWidth-1: AddrWidth-ReminderBits];
    assign aw_const    = dram_req_interleaved[i].aw.addr[ConstantBits-1 : 0];

    if (NumDrams == 1) begin
      assign aw_scramble_addr_reset = {aw_reminder, aw_scramble, aw_const};
    end else begin
      assign aw_scramble_addr_reset = {{ScrambleBits{1'b0}}, aw_reminder, aw_const};
    end

    // req.ar scrambling
    logic [ConstantBits-1:0] ar_const;
    logic [ScrambleBits-1:0] ar_scramble;
    logic [ReminderBits-1:0] ar_reminder;
    logic [AddrWidth-1   :0] ar_scramble_addr_reset;
    assign ar_scramble = dram_req_interleaved[i].ar.addr[AddrWidth-1 : AddrWidth-ScrambleBits];
    assign ar_reminder = dram_req_interleaved[i].ar.addr[AddrWidth-ScrambleBits-1 : ConstantBits] - L2MemoryBaseAddr[AddrWidth-1: AddrWidth-ReminderBits];
    assign ar_const    = dram_req_interleaved[i].ar.addr[ConstantBits-1 : 0];

    if (NumDrams == 1) begin
      assign ar_scramble_addr_reset = {ar_reminder, ar_scramble, ar_const};
    end else begin
      assign ar_scramble_addr_reset = {{ScrambleBits{1'b0}}, ar_reminder, ar_const};
    end

    // Scrambled AXI req assignment
    always_comb begin
      dram_req[i]         = dram_req_interleaved[i];
      dram_req[i].aw.addr = aw_scramble_addr_reset;
      dram_req[i].ar.addr = ar_scramble_addr_reset;
    end
  end: gen_dram_scrambler_reset

  for (genvar i = 0; unsigned'(i) < NumDrams; i++) begin: gen_drams
    axi_dram_sim #(
        .AxiAddrWidth(AddrWidth        ),
        .AxiDataWidth(AxiDataWidth     ),
        .AxiIdWidth  (AxiSystemIdWidth ),
        .AxiUserWidth(1                ),
        .BASE        ('b0              ),
        .axi_req_t   (axi_system_req_t ),
        .axi_resp_t  (axi_system_resp_t),
        .axi_ar_t    (axi_system_ar_t  ),
        .axi_r_t     (axi_system_r_t   ),
        .axi_aw_t    (axi_system_aw_t  ),
        .axi_w_t     (axi_system_w_t   ),
        .axi_b_t     (axi_system_b_t   )
    ) i_axi_dram_sim (
        .clk_i,
        .rst_ni,
        .axi_req_i (dram_req[i] ),
        .axi_resp_o(dram_resp[i])
    );
  end: gen_drams
`endif

  /*************
   *  Bootrom  *
   *************/

  // Memory
  logic      bootrom_req;
  logic      bootrom_rvalid;
  addr_t     bootrom_addr;
  axi_data_t bootrom_rdata;

  axi2mem #(
    .axi_req_t  (axi_system_req_t ),
    .axi_resp_t (axi_system_resp_t),
    .AddrWidth  (AddrWidth        ),
    .DataWidth  (AxiDataWidth     ),
    .IdWidth    (AxiSystemIdWidth ),
    .NumBanks   (1                ),
    .BufDepth   (2                )
  ) i_axi2mem_bootrom (
    .clk_i        (clk_i                   ),
    .rst_ni       (rst_ni                  ),

    .busy_o       (/*unsused*/             ),

    .axi_req_i    (axi_periph_req[Bootrom] ),
    .axi_resp_o   (axi_periph_resp[Bootrom]),

    .mem_req_o    (bootrom_req             ),
    .mem_gnt_i    (bootrom_req             ),
    .mem_addr_o   (bootrom_addr            ),
    .mem_wdata_o  (/*unused*/              ),
    .mem_strb_o   (/*unused*/              ),
    .mem_atop_o   (/*unused*/              ),
    .mem_we_o     (/*unused*/              ),
    .mem_rvalid_i (bootrom_rvalid          ),
    .mem_rdata_i  (bootrom_rdata           )
  );

  `FF(bootrom_rvalid, bootrom_req, 1'b0, clk_i, rst_ni)

  bootrom i_bootrom (
    .clk_i  (clk_i        ),
    .req_i  (bootrom_req  ),
    .addr_i (bootrom_addr ),
    .rdata_o(bootrom_rdata)
  );

  /***********************
   *  Control Registers  *
   ***********************/

  localparam NumPeriphs = 2; // Control registers + DMA

  typedef enum logic [$clog2(NumPeriphs) - 1:0] {
    CtrlRegisters,
    DMA
  } axi_lite_xbar_slave_target;

  axi_periph_req_t                     axi_periph_narrow_req;
  axi_periph_resp_t                    axi_periph_narrow_resp;
  axi_periph_req_t    [NumClusters-1:0] axi_demuxed_narrow_req;
  axi_periph_resp_t   [NumClusters-1:0] axi_demuxed_narrow_resp;
  axi_lite_slv_req_t  [NumClusters-1:0] axi_lite_mst_req;
  axi_lite_slv_resp_t [NumClusters-1:0] axi_lite_mst_resp;
  axi_lite_slv_req_t  [NumClusters-1:0][NumPeriphs-1:0] axi_lite_slv_req;
  axi_lite_slv_resp_t [NumClusters-1:0][NumPeriphs-1:0] axi_lite_slv_resp;



  localparam xbar_cfg_t AXILiteXBarCfg = '{
    NoSlvPorts         : 1,
    NoMstPorts         : NumPeriphs,
    MaxMstTrans        : 1,
    MaxSlvTrans        : 1,
    FallThrough        : 1'b0,
    LatencyMode        : axi_pkg::NO_LATENCY,
    PipelineStages     : 0,
    AxiIdWidthSlvPorts : 0, /* Not used for AXI lite */
    AxiIdUsedSlvPorts  : 0, /* Not used for AXI lite */
    UniqueIds          : 0, /* Not used for AXI lite */
    AxiAddrWidth       : AddrWidth,
    AxiDataWidth       : AxiLiteDataWidth,
    NoAddrRules        : NumPeriphs
  };

  localparam addr_t CtrlRegistersBaseAddr = 32'h4000_0000;
  localparam addr_t CtrlRegistersEndAddr  = 32'h4001_0000;
  localparam addr_t DMABaseAddr           = 32'h4001_0000;
  localparam addr_t DMAEndAddr            = 32'h4002_0000;

  xbar_rule_32_t [NumPeriphs-1:0] axi_lite_xbar_rules;
  assign axi_lite_xbar_rules = '{
    '{idx: CtrlRegisters, start_addr: CtrlRegistersBaseAddr, end_addr: CtrlRegistersEndAddr},
    '{idx: DMA, start_addr: DMABaseAddr, end_addr: DMAEndAddr}
  };

  axi_dw_converter #(
    .AxiMaxReads         (1                ), // Number of outstanding reads
    .AxiSlvPortDataWidth (AxiDataWidth     ), // Data width of the slv port
    .AxiMstPortDataWidth (AxiLiteDataWidth ), // Data width of the mst port
    .AxiAddrWidth        (AddrWidth        ), // Address width
    .AxiIdWidth          (AxiSystemIdWidth ), // ID width
    .aw_chan_t           (axi_system_aw_t  ), // AW Channel Type
    .mst_w_chan_t        (axi_periph_w_t   ), //  W Channel Type for the mst port
    .slv_w_chan_t        (axi_system_w_t   ), //  W Channel Type for the slv port
    .b_chan_t            (axi_system_b_t   ), //  B Channel Type
    .ar_chan_t           (axi_system_ar_t  ), // AR Channel Type
    .mst_r_chan_t        (axi_periph_r_t   ), //  R Channel Type for the mst port
    .slv_r_chan_t        (axi_system_r_t   ), //  R Channel Type for the slv port
    .axi_mst_req_t       (axi_periph_req_t ), // AXI Request Type for mst ports
    .axi_mst_resp_t      (axi_periph_resp_t), // AXI Response Type for mst ports
    .axi_slv_req_t       (axi_system_req_t ), // AXI Request Type for slv ports
    .axi_slv_resp_t      (axi_system_resp_t)  // AXI Response Type for slv ports
  ) i_axi_dw_converter_ctrl (
    .clk_i      (clk_i                       ),
    .rst_ni     (rst_ni                      ),
    // Slave interface
    .slv_req_i  (axi_periph_req[Peripherals] ),
    .slv_resp_o (axi_periph_resp[Peripherals]),
    // Master interface
    .mst_req_o  (axi_periph_narrow_req       ),
    .mst_resp_i (axi_periph_narrow_resp      )
  );

  // Demux AXI signal between peripherals for each cluster
  axi_demux #(
    .AxiIdWidth          (AxiSystemIdWidth ), // ID width
    .aw_chan_t           (axi_system_aw_t  ), // AW Channel Type
    .w_chan_t            (axi_periph_w_t   ), //  W Channel Type
    .b_chan_t            (axi_system_b_t   ), //  B Channel Type
    .ar_chan_t           (axi_system_ar_t  ), // AR Channel Type
    .r_chan_t            (axi_periph_r_t   ), //  R Channel Type
    .axi_req_t           (axi_periph_req_t ), // AXI Request Type
    .axi_resp_t          (axi_periph_resp_t), // AXI Response Type
    .NoMstPorts (NumClusters        ), // Number of instantiated ports
    .MaxTrans   (4                  )  // Maximum number of open transactions per channel
  ) axi_periph_demux_i(
    .clk_i            (clk_i                         ),
    .rst_ni           (rst_ni                        ),
    .test_i           (/*unused*/                    ),
    // Slave Port
    .slv_req_i        (axi_periph_narrow_req         ),
    .slv_aw_select_i  (axi_periph_narrow_req.aw.user  ),
    .slv_ar_select_i  (axi_periph_narrow_req.ar.user ),
    .slv_resp_o       (axi_periph_narrow_resp        ),
    // Master Ports
    .mst_reqs_o       (axi_demuxed_narrow_req        ),
    .mst_resps_i      (axi_demuxed_narrow_resp       )
  );

  // Generate cluster peripherals
  for(genvar i = 0; i < NumClusters; i++) begin: gen_cluster_peripherals

    axi_to_axi_lite #(
      .AxiAddrWidth   (AddrWidth          ),
      .AxiDataWidth   (AxiLiteDataWidth   ),
      .AxiIdWidth     (AxiSystemIdWidth   ),
      .AxiUserWidth   (1                  ),
      .AxiMaxReadTxns (1                  ),
      .AxiMaxWriteTxns(1                  ),
      .FallThrough    (1'b0               ),
      .full_req_t     (axi_periph_req_t   ),
      .full_resp_t    (axi_periph_resp_t  ),
      .lite_req_t     (axi_lite_slv_req_t ),
      .lite_resp_t    (axi_lite_slv_resp_t)
    ) i_axi_to_axi_lite (
      .clk_i     (clk_i                     ),
      .rst_ni    (rst_ni                    ),
      .test_i    (1'b0                      ),
      .slv_req_i (axi_demuxed_narrow_req[i] ),
      .slv_resp_o(axi_demuxed_narrow_resp[i]),
      .mst_req_o (axi_lite_mst_req[i]       ),
      .mst_resp_i(axi_lite_mst_resp[i]      )
    );
    axi_lite_xbar #(
      .Cfg       (AXILiteXBarCfg     ),
      .aw_chan_t (axi_lite_slv_aw_t  ),
      .w_chan_t  (axi_lite_slv_w_t   ),
      .b_chan_t  (axi_lite_slv_b_t   ),
      .ar_chan_t (axi_lite_slv_ar_t  ),
      .r_chan_t  (axi_lite_slv_r_t   ),
      .axi_req_t (axi_lite_slv_req_t ),
      .axi_resp_t(axi_lite_slv_resp_t),
      .rule_t    (xbar_rule_32_t     )
    ) i_axi_lite_xbar (
      .clk_i                (clk_i                 ),
      .rst_ni               (rst_ni                ),
      .test_i               (1'b0                  ),
      .slv_ports_req_i      (axi_lite_mst_req[i]   ),
      .slv_ports_resp_o     (axi_lite_mst_resp[i]  ),
      .mst_ports_req_o      (axi_lite_slv_req[i]   ),
      .mst_ports_resp_i     (axi_lite_slv_resp[i]  ),
      .addr_map_i           (axi_lite_xbar_rules   ),
      .en_default_mst_port_i('1                    ),
      .default_mst_port_i   (CtrlRegisters         )
    );

    ctrl_registers #(
      .NumRegs          (16 + 8             ),
      .TCDMBaseAddr     (TCDMBaseAddr       ),
      .TCDMSize         (TCDMSize           ),
      .NumCores         (NumCores           ),
      .axi_lite_req_t (axi_lite_slv_req_t ),
      .axi_lite_resp_t(axi_lite_slv_resp_t)
    ) i_ctrl_registers (
      .clk_i                (clk_i                               ),
      .rst_ni               (rst_ni                              ),
      .axi_lite_slave_req_i (axi_lite_slv_req[i][CtrlRegisters]  ),
      .axi_lite_slave_resp_o(axi_lite_slv_resp[i][CtrlRegisters] ),
      .ro_cache_ctrl_o      (ro_cache_ctrl[i]                    ),
      .tcdm_start_address_o (/* Unused */                        ),
      .tcdm_end_address_o   (/* Unused */                        ),
      .num_cores_o          (/* Unused */                        ),
      .wake_up_o            (wake_up[i]                          ),
      .eoc_o                (/* Unused */                        ),
      .eoc_valid_o          (eoc_valid[i]                        )
    );
    mempool_dma #(
      .axi_lite_req_t(axi_lite_slv_req_t       ),
      .axi_lite_rsp_t(axi_lite_slv_resp_t      ),
      .burst_req_t   (dma_req_t                ),
      .NumBackends   (NumGroups                ),
      .DmaIdWidth    (1                        )
    ) i_mempool_dma (
      .clk_i           (clk_i                           ),
      .rst_ni          (rst_ni                          ),
      .config_req_i    (axi_lite_slv_req[i][DMA]        ),
      .config_res_o    (axi_lite_slv_resp[i][DMA]       ),
      .burst_req_o     (dma_req[i]                      ),
      .valid_o         (dma_req_valid[i]                ),
      .ready_i         (dma_req_ready[i]                ),
      .backend_idle_i  (dma_meta[i].backend_idle        ),
      .trans_complete_i(dma_meta[i].trans_complete      ),
      .dma_id_o        (dma_id[i]                       )
    );
  end

  assign busy_o = 1'b0;

  // From MemPool to the Host
  assign mst_req_o                 = axi_periph_req[External];
  assign axi_periph_resp[External] = mst_resp_i;
  // From the Host to MemPool
  axi_id_remap #(
    .AxiSlvPortIdWidth   (AxiSystemIdWidth ),
    .AxiSlvPortMaxUniqIds(1                ),
    .AxiMaxTxnsPerId     (1                ),
    .AxiMstPortIdWidth   (AxiTileIdWidth   ),
    .slv_req_t           (axi_system_req_t ),
    .slv_resp_t          (axi_system_resp_t),
    .mst_req_t           (axi_tile_req_t   ),
    .mst_resp_t          (axi_tile_resp_t  )
  ) i_axi_id_remap (
    .clk_i     (clk_i                        ),
    .rst_ni    (rst_ni                       ),
    .slv_req_i (slv_req_i                    ),
    .slv_resp_o(slv_resp_o                   ),
    .mst_req_o (axi_mst_req[NumSystemXbarMasters-1] ),
    .mst_resp_i(axi_mst_resp[NumSystemXbarMasters-1])
  );

endmodule : mempool_system
