../../../../toolchain/riscv-opcodes/inst.sverilog