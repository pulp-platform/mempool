../../tb_tcdm_interconnect/hdl/defaults.svh