../riscv-opcodes/inst.sverilog