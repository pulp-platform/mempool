../../tb_tcdm_interconnect/hdl/tb_patterns.sv